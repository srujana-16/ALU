`timescale 1ns / 1ps

module xor_TB;


reg signed[63:0] a,b;
wire signed[63:0] y;

bitxor uut(
    .a(a),
    .b(b),
    .y(y)
);

initial begin 
		$dumpfile("bitxor.vcd");
     	$dumpvars(0,xor_TB);
		
    a = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    b = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    #100;
    a = 64'b0000000000000000000000000000000000000000000000000000010000000101;
    b = 64'b0000000000000000000000000000000000000000000000000000010000000011;
    #20;
    a = 64'b0000000000000000000000000000000000000000000000000101110110011111;
    b = 64'b0000000000000000000000000000000000000000000011110000110010110010;
    #20;
    a = 64'b0000000000000000000000000000000000000000000000000010010000110101;
    b = 64'b1111111111111111111100001000100000000000000000000000000000000000;
    #20;
    a = 64'b1111111111110011111001110011111100000000000000000000000000000000;
    b = 64'b0000000000000000000010101011011100000000000000000000000000000000;
    #20;
    a = 64'b1111111111110011110000000011100000000000000000000000000000000000;
    b = 64'b1111111111111111111101111110110100000000000000000000000000000000;
    #20;

     
end 
    initial begin 
        $monitor("a=%d b=%d y=%d\n",a,b,y);
        end 

endmodule