`timescale 1ns / 1ps

module ALU_TB;

reg [1:0] Control;
reg signed [63:0] a,b;
wire signed [63:0] y;

ALU uut(
    .Control(Control),
    .a(a),
    .b(b),
    .y(y)
);

initial begin 
		$dumpfile("ALU.vcd");
     	$dumpvars(0,ALU_TB);
	
    a=0;
    b=0;
    Control=0;	
    #100; 
    a = 64'b0000000000000000000000000000000000000000000000000000010000000101;
    b = 64'b0000000000000000000000000000000000000000000000000000010000000011;
    Control = 2'b00; 
    #20 Control = 2'b01;
    #20 Control = 2'b10;
    #20 Control = 2'b11;
    #20;
    a = 64'b0000000000000000000000000000000000000000000000000101110110011111;
    b = 64'b0000000000000000000000000000000000000000000011110000110010110010;
    Control = 2'b00; 
    #20 Control = 2'b01;
    #20 Control = 2'b10;
    #20 Control = 2'b11;
    #20;
    a = 64'b0000000000000000000000000000000000000000000000000010010000110101;
    b = 64'b1111111111111111111100001000100000000000000000000000000000000000;
    Control = 2'b00; 
    #20 Control = 2'b01;
    #20 Control = 2'b10;
    #20 Control = 2'b11;
    #20;
    a = 64'b1111111111110011111001110011111100000000000000000000000000000000;
    b = 64'b0000000000000000000010101011011100000000000000000000000000000000;
    Control = 2'b00; 
    #20 Control = 2'b01;
    #20 Control = 2'b10;
    #20 Control = 2'b11;
    #20;
    a = 64'b1111111111110011110000000011100000000000000000000000000000000000;
    b = 64'b1111111111111111111101111110110100000000000000000000000000000000;
    Control = 2'b00; 
    #20 Control = 2'b01;
    #20 Control = 2'b10;
    #20 Control = 2'b11;
    #20;
    end
      initial begin 
        $monitor("a=%d b=%d Control=%d y=%d\n",a,b,Control,y);
        end 

endmodule